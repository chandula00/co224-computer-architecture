// Computer Architecture (CO224) - Lab 05
// Design: Testbench of Integrated CPU of Simple Processor
// Author: Isuru Nawinne

// simulation time will advance by 1 nanosecond for every 100 picoseconds of real time
`timescale 1ns/100ps

`include "cpu.v"
`include "dmem.v"
`include "dcache.v"
`include "imem.v"
`include "icache.v"

module cpu_tb;

    reg CLK, RESET;
    wire [31:0] PC;
    wire [31:0] INSTRUCTION;
    
    
    wire CPU_READ, CPU_WRITE, CPU_BUSYWAIT;
	wire DM_READ, DM_WRITE, DM_BUSYWAIT, DC_BUSYWAIT;
    wire IM_READ, IM_BUSYWAIT, IC_BUSYWAIT;
	
	wire [7:0] CPU_ADDRESS, CPU_WRITEDATA, CPU_READDATA;
	wire [31:0] DM_WRITEDATA, DM_READDATA;
	wire [5:0] DM_ADDRESS;
    
    wire [5:0] IM_ADDRESS;
	wire [127:0] IM_INSTR;
    /* 
    ------------------------
     SIMPLE INSTRUCTION MEM
    ------------------------
    */
    
    // // TODO: Initialize an array of registers (8x1024) named 'instr_mem' to be used as instruction memory
    // reg [7:0] instr_mem [1023:0];
    
    // // TODO: Create combinational logic to support CPU instruction fetching, given the Program Counter(PC) value 
    // //       (make sure you include the delay for instruction fetching here)
    // assign #2 INSTRUCTION = {instr_mem[PC+3],instr_mem[PC+2],instr_mem[PC+1],instr_mem[PC]};
    
    // initial
    // begin
    //     // Initialize instruction memory with the set of instructions you need execute on CPU
        
    //     // METHOD 1: manually loading instructions to instr_mem
    //     //{instr_mem[10'd3], instr_mem[10'd2], instr_mem[10'd1], instr_mem[10'd0]} = 32'b00000000000001000000000000000101;
    //     //{instr_mem[10'd7], instr_mem[10'd6], instr_mem[10'd5], instr_mem[10'd4]} = 32'b00000000000000100000000000001001;
    //     //{instr_mem[10'd11], instr_mem[10'd10], instr_mem[10'd9], instr_mem[10'd8]} = 32'b00000010000001100000010000000010;
        
    //     // METHOD 2: loading instr_mem content from instr_mem.mem file
    //     $readmemb("instr_mem.mem", instr_mem);
    //     //$display("instr_mem = %h",instr_mem);
    // end
    
    
    /*
	------------
	DATA MEMORY
	------------
    */
	dataMemory mydatamem(CLK, RESET, DM_READ, DM_WRITE, DM_ADDRESS, DM_WRITEDATA, DM_READDATA, DM_BUSYWAIT);
	
	/*
	------------
	DATA CACHE
	------------
    */
	dcache mydatacache (CLK, RESET, CPU_READ, CPU_WRITE, CPU_ADDRESS, CPU_WRITEDATA, CPU_READDATA, DC_BUSYWAIT, DM_READ, DM_WRITE, DM_ADDRESS, DM_WRITEDATA, DM_READDATA, DM_BUSYWAIT);

    /*
	------------------
	INSTRUCTION CACHE
	------------------
    */
	icache myicache(CLK, RESET, PC[9:0], INSTRUCTION, IC_BUSYWAIT, IM_READ, IM_ADDRESS, IM_INSTR, IM_BUSYWAIT);
	
	/*
	------------------
	INSTRUCTION MEMORY
	------------------
    */
	imemory myimemory(CLK, IM_READ, IM_ADDRESS, IM_INSTR, IM_BUSYWAIT);
    assign CPU_BUSYWAIT = IC_BUSYWAIT || DC_BUSYWAIT;
    /* 
    -----
     CPU
    -----
    */
    cpu mycpu(PC, INSTRUCTION, CLK, RESET, CPU_READ, CPU_WRITE, CPU_ADDRESS, CPU_WRITEDATA, CPU_READDATA, CPU_BUSYWAIT);

    initial
    begin
    
        // generate files needed to plot the waveform using GTKWave
        $dumpfile("cpu_wavedata.vcd");
		$dumpvars(0, cpu_tb);
        
        CLK = 1'b0;
        RESET = 1'b0;
        
        // TODO: Reset the CPU (by giving a pulse to RESET signal) to start the program execution
        RESET = 1'b1;
		#5
		RESET = 1'b0;


        // finish simulation after some time
        #5000
        $finish;
        
    end
    
    // clock signal generation
    always
        #4 CLK = ~CLK;
        

endmodule